module main
const (
    icons = {
        "git_branch": "\ue725"
        "git_ahead": "\ufc35",
        "git_staged": "\uf42e",
        "git_unstaged": "\uf8ea",
        "git_untracked": "\uf44d",
        "git_conflicted": "\ue727",
        "git_stash": "\uf187"
    }
)
