
module main

const (
	init_bg = 237
	init_fg = 254 
	user_bg = 153
	user_fg = 238

	cmd_s_bg = 40
	cmd_s_fg = 238
	cmd_f_bg = 161
	cmd_f_fg = 238

	cwd_bg = 237
	cwd_fg = 254 

	git_master_bg = 206
	git_branch_bg = 153
	git_branch_fg = 238
)