
module main

const (
    init_bg = 237
    init_fg = 254 
    user_bg = 153
    user_fg = 238

    cmd_s_bg = 77
    cmd_s_fg = 238
    cmd_f_bg = 126
    cmd_f_fg = 238

    cwd_bg = 237
    cwd_fg = 254 

    git_master_bg = 75
    git_branch_bg = 65
    git_branch_fg = 238

    staged_bg = 120
    staged_fg = 238
    unstaged_bg = 213
    unstaged_fg = 238
    untracked_bg = 88
    untracked_fg = 255
)
