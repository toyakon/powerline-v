
module main

const (
	user_bg = 153
	user_fg = 238

	cmd_s_bg = 153
	cmd_s_fg = 238
	cmd_f_bg = 161
	cmd_f_fg = 238
)